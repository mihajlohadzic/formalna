bind zadaci a_checker c0(.clk(clk), .rst(rst), .rt(rt), .rdy(rdy), .start(start), .endd(endd)
, .er2(er2), .er3(er3), .rdy3(rdy3), .rdy4(rdy4), .start4(start4), .endd5(endd5), .stop5(stop5),
.er5(er5), .rdy5(rdy5), .start5(start5), .endd6(endd6), .stop6(stop6),.er6(er6),.rdy6(rdy6),.endd7(endd7),
.start7(start7),.status_valid7(status_valid7),.instartsv7(instartsv7),.rt8(rt8),.enable8(enable8),.rdy9(rdy9),.start9(start9),
.interrupt9(interrupt9), .ack10(ack10), .req10(req10)
);