bind zadaci a_checker c0(.clk(clk), .rst(rst), .rt(rt), .rdy(rdy), .start(start), .endd(endd)
, .er2(er2), .er3(er3), .rdy3(rdy3), .rdy4(rdy4), .start4(start4), .endd5(endd5), .stop5(stop5),
.er5(er5), .rdy5(rdy5), .start5(start5)
);